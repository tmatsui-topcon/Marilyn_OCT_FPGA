-- ***************************************************************************************
--		******  Copyright (c) 2007 by TOPCON Corp.  All rights reserved.  ******		--
-- ***************************************************************************************
-- File name			:H_W_Rev.vhd : VHDL File
-- Detail of Function	:FPGAハードウェアレビジョン通知回路
-- Date					:070808
-- Created by			:Y.NISHIO
--<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<< Change history >>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>
-- [2007/08/08 : H_W_Rev_001]
--  ・新規作成
-- [2007/10/12]
--  ・ハードウェアバージョンの設定値入力を16進に変更
--
--
-- [2018/03/16]ver1.0.0.2
--  ・ガルバノ波形乱れ対応
--    MaetstroのOCT基板FPGAver1.1.1.3で対応された内容を反映 T.Sato
--
--**************************************************************************************--
--********************	Library declaration part			****************************--
--**************************************************************************************--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

--**************************************************************************************--
--********************	Entity Declaration					****************************--
--**************************************************************************************--
entity H_W_Rev is
	port(
		H_W_Rev_1	:	out	std_logic_vector(3 downto 0);
		H_W_Rev_2	:	out	std_logic_vector(3 downto 0);
		H_W_Rev_3	:	out	std_logic_vector(3 downto 0);
		H_W_Rev_4	:	out	std_logic_vector(3 downto 0)
	);
end H_W_Rev;

--**************************************************************************************--
--********************	Architecture Body					****************************--
--**************************************************************************************--
architecture RTL of H_W_Rev is

--**************************************************************************************--
--********************	Signal definition part				****************************--
--**************************************************************************************--
	constant	const_H_W_Rev_1:	std_logic_vector(3 downto 0) := X"0";
	constant	const_H_W_Rev_2:	std_logic_vector(3 downto 0) := X"0";
	constant	const_H_W_Rev_3:	std_logic_vector(3 downto 0) := X"0";
	constant	const_H_W_Rev_4:	std_logic_vector(3 downto 0) := X"9";

--**************************************************************************************--
begin

--*************** ハードウェアバージョン出力 ******************************************--
	H_W_Rev_1	<= const_H_W_Rev_1;
	H_W_Rev_2	<= const_H_W_Rev_2;
	H_W_Rev_3	<= const_H_W_Rev_3;
	H_W_Rev_4	<= const_H_W_Rev_4;
-----------------------------------------------------------------------------------------
end RTL;
