-- ***************************************************************************************
--		******  Copyright (c) 2007 by TOPCON Corp.  All rights reserved.  ******		--
-- ***************************************************************************************
-- File name			:comp_TRIG_SEL.vhd : VHDL File			-- <<<<<< Check Version
-- Ver					:001									-- <<<<<< Check Version
-- Date					:20081104
-- Created by			:�k�h�s�Z�l����
--<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<< Change history >>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>
-- [2008/11/04 : comp_TRIG_001]
--	1.TRIG�I�����W���[��
--		�J�X�^���X�L�����p�R���|�[�l���g
--
--
--**************************************************************************************--
--********************	Library declaration part			****************************--
--**************************************************************************************--
LIBRARY ieee;
LIBRARY lpm;
LIBRARY altera_mf;
USE ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

--**************************************************************************************--
--********************	Entity Declaration					****************************--
--**************************************************************************************--
ENTITY comp_TRIG_SEL IS
	PORT
	(
		FPGAclk : IN STD_LOGIC;						--20MHz
		Reset : IN STD_LOGIC;
		TRIG_IN :  IN STD_LOGIC;	--from galv_con
		TRIG_EN : IN STD_LOGIC;
		Custom_Flag : IN STD_LOGIC;
		TRIG_OUT : OUT STD_LOGIC
		);
END  comp_TRIG_SEL;

--**************************************************************************************--
--********************	Architecture Body					****************************--
--**************************************************************************************--
ARCHITECTURE RTL OF comp_TRIG_SEL IS

--**************************************************************************************--
--********************	Signal definition part				****************************--
--**************************************************************************************--
	signal sig_TRIG_OUT : std_logic;

-----------------------------------------------------------------------------------------
begin

-----------------------------------------------------------------------------------------
	TRIG_OUT <= sig_TRIG_OUT;

-----------------------------------------------------------------------------------------
	U_TRIG_OUT :
	process(
		Reset,
		FPGAclk
	) begin
		if(
			Reset = '1'
		) then
			sig_TRIG_OUT <= '0';
		elsif(
			FPGAclk'event and FPGAclk='1'
		) then
			if(
				Custom_Flag = '0'
			) then
				sig_TRIG_OUT <= TRIG_IN;
			else
				if(
					TRIG_EN = '1'
				) then
					if( TRIG_IN = '1' )then
						sig_TRIG_OUT <= '1';
					end if;
				else
					sig_TRIG_OUT <= '0';
				end if;
			end if;
		end if;
	end process;

-----------------------------------------------------------------------------------------
END RTL;
