-- ***************************************************************************************
--		******  Copyright (c) 2015 by TOPCON Corp.  All rights reserved.  ******		--
-- ***************************************************************************************
--
--
--**************************************************************************************--
--********************	Library declaration part			****************************--
--**************************************************************************************--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

--**************************************************************************************--
--********************	Entity Declaration					****************************--
--**************************************************************************************--
entity make_abs is
	port(
		FPGAclk		:	in	std_logic;
		Reset		:	in	std_logic;
		data_i		:	in	std_logic_vector(15 downto 0);
		data_o		:	out	std_logic_vector(15 downto 0)
	);
end make_abs;

--**************************************************************************************--
--********************	Architecture Body					****************************--
--**************************************************************************************--
architecture RTL of make_abs is


--**************************************************************************************--
--********************	Signal definition part				****************************--
--**************************************************************************************--
	signal	reg_abs_data		: std_logic_vector(15 downto 0);

begin
	data_o <= reg_abs_data;

	process( Reset, FPGAclk) 
	begin
		if( Reset = '1') then
			reg_abs_data <= (others => '0');
		elsif( FPGAclk'event and FPGAclk='1') then
			if(data_i(15) = '1')then
				reg_abs_data <= not data_i + X"0001";
			else
				reg_abs_data <= data_i ;
			end if;
		end if;
	end process;
	
-----------------------------------------------------------------------------------------
end RTL;
